library verilog;
use verilog.vl_types.all;
entity Peaje_vlg_vec_tst is
end Peaje_vlg_vec_tst;

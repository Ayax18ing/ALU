library verilog;
use verilog.vl_types.all;
entity Sem_fin_vlg_check_tst is
    port(
        rojo            : in     vl_logic;
        talfin          : in     vl_logic;
        verde           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Sem_fin_vlg_check_tst;

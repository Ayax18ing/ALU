library verilog;
use verilog.vl_types.all;
entity Back_sensor_vlg_vec_tst is
end Back_sensor_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity contador_vehiculos_vlg_vec_tst is
end contador_vehiculos_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Parcial_2_vlg_vec_tst is
end Parcial_2_vlg_vec_tst;

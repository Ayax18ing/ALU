library verilog;
use verilog.vl_types.all;
entity Contador_as_vlg_vec_tst is
end Contador_as_vlg_vec_tst;

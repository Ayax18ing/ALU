library verilog;
use verilog.vl_types.all;
entity Sem_fin_vlg_vec_tst is
end Sem_fin_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity ALU_E_vlg_vec_tst is
end ALU_E_vlg_vec_tst;

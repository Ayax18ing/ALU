library verilog;
use verilog.vl_types.all;
entity Contador_tiempo_vlg_vec_tst is
end Contador_tiempo_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Front_sensor_vlg_vec_tst is
end Front_sensor_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Contador_des_vlg_vec_tst is
end Contador_des_vlg_vec_tst;
